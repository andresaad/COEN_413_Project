library verilog;
use verilog.vl_types.all;
entity root_sv_unit is
end root_sv_unit;
