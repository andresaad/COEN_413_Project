library verilog;
use verilog.vl_types.all;
entity test_02_constrained_sv_unit is
end test_02_constrained_sv_unit;
