library verilog;
use verilog.vl_types.all;
entity calc2_if is
    port(
        PClk            : in     vl_logic
    );
end calc2_if;
