parameter CALC_CMD_WIDTH = 4;
typedef bit [CALC_CMD_WIDTH-1:0] reg_cmd_t;
parameter CALC_DATA_WIDTH = 32;
typedef bit [CALC_DATA_WIDTH-1:0] req_data_t;
