library verilog;
use verilog.vl_types.all;
entity scoreboard_sv_unit is
end scoreboard_sv_unit;
