library verilog;
use verilog.vl_types.all;
entity test_03_cvr_driven_sv_unit is
end test_03_cvr_driven_sv_unit;
