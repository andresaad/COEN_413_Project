library verilog;
use verilog.vl_types.all;
entity test_01_directed_sv_unit is
end test_01_directed_sv_unit;
