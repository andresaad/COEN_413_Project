library verilog;
use verilog.vl_types.all;
entity apb_if_sv_unit is
end apb_if_sv_unit;
