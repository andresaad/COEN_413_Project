library verilog;
use verilog.vl_types.all;
entity apb_if is
    port(
        PClk            : in     vl_logic
    );
end apb_if;
