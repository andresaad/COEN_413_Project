library verilog;
use verilog.vl_types.all;
entity apb_trans_sv_unit is
end apb_trans_sv_unit;
