library verilog;
use verilog.vl_types.all;
entity calc_result_sv_unit is
end calc_result_sv_unit;
