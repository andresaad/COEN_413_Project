library verilog;
use verilog.vl_types.all;
entity calc_master_sv_unit is
end calc_master_sv_unit;
