library verilog;
use verilog.vl_types.all;
entity request_gen_sv_unit is
end request_gen_sv_unit;
