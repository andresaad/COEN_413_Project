library verilog;
use verilog.vl_types.all;
entity apb_gen_sv_unit is
end apb_gen_sv_unit;
