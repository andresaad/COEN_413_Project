// Root File, Stores data and adresse width

parameter APB_ADDR_WIDTH = 16;
typedef bit [APB_ADDR_WIDTH-1:0] apb_addr_t;
parameter APB_WIDTH = 32;
typedef bit [APB_WIDTH-1:0] app_data_t;
typedef enum {READ, WRITE, IDLE} transe_e;
