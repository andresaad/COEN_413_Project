library verilog;
use verilog.vl_types.all;
entity apb_monitor_sv_unit is
end apb_monitor_sv_unit;
