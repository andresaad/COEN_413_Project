library verilog;
use verilog.vl_types.all;
entity testbench_sv_unit is
end testbench_sv_unit;
