library verilog;
use verilog.vl_types.all;
entity apb_result_sv_unit is
end apb_result_sv_unit;
