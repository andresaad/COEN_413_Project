library verilog;
use verilog.vl_types.all;
entity apb_master_sv_unit is
end apb_master_sv_unit;
