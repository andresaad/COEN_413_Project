library verilog;
use verilog.vl_types.all;
entity Master_sv_unit is
end Master_sv_unit;
