library verilog;
use verilog.vl_types.all;
entity Rslt_sv_unit is
end Rslt_sv_unit;
