library verilog;
use verilog.vl_types.all;
entity calc2_if_sv_unit is
end calc2_if_sv_unit;
