library verilog;
use verilog.vl_types.all;
entity calc_monitor_sv_unit is
end calc_monitor_sv_unit;
