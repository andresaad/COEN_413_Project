library verilog;
use verilog.vl_types.all;
entity mem_sv_unit is
end mem_sv_unit;
