library verilog;
use verilog.vl_types.all;
entity mem is
end mem;
