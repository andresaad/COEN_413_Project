library verilog;
use verilog.vl_types.all;
entity calc_request_sv_unit is
end calc_request_sv_unit;
